module decoder1_2(input d,output y0,y1);
  assign y0 = ~d;
  assign y1 = d;
endmodule
