module mux4_1_tb;
  reg i0,i1,i2,i3,s0,s1;
  wire y;
  mux4_1 dut(.*);
  initial begin
    $dumpfile("mux4_1.vcd");
    $dumpvars(1,mux4_1_tb);
    $monitor("$time=0%t i0=%b i1=%b i2=%b i3=%b s0=%b s1=%b y=%b",$time,i0,i1,i2,i3,s0,s1,y);
    i0=1; i1=0; i2=1; i3=0;
    s0=0; s1=0; #10
    s0=0; s1=1; #10
    s0=1; s1=0; #10
    s0=1; s1=1; #10
    $finish;
  end
endmodule
    
    
