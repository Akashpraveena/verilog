module demux1_4(input din,input [1:0]s , output reg y0,y1,y2,y3);
  always@(*) begin
    y0 = 0;
    y1 = 0;
    y2 = 0;
    y3 = 0;
     case(s)
       2'b00 : y0 = din;
       2'b01 : y1 = din;
       2'b10 : y2 = din;
       2'b11 : y3 = din;
    endcase
  end 
endmodule
      
